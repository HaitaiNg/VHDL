

# PlanAhead Generated physical constraints

NET "an[7]" LOC = U13;
NET "an[6]" LOC = K2;
NET "an[5]" LOC = T14;
NET "an[4]" LOC = P14;
NET "an[3]" LOC = J14;
NET "an[2]" LOC = T9;
NET "an[1]" LOC = J18;
NET "an[0]" LOC = J17;

# PlanAhead Generated IO constraints

NET "an[7]" IOSTANDARD = LVCMOS33;
NET "an[6]" IOSTANDARD = LVCMOS33;
NET "an[5]" IOSTANDARD = LVCMOS33;
NET "an[4]" IOSTANDARD = LVCMOS33;
NET "an[3]" IOSTANDARD = LVCMOS33;
NET "an[2]" IOSTANDARD = LVCMOS33;
NET "an[1]" IOSTANDARD = LVCMOS33;
NET "an[0]" IOSTANDARD = LVCMOS33;
NET "sseg_sign[6]" IOSTANDARD = LVCMOS33;
NET "sseg_sign[5]" IOSTANDARD = LVCMOS33;
NET "sseg_sign[4]" IOSTANDARD = LVCMOS33;
NET "sseg_sign[3]" IOSTANDARD = LVCMOS33;
NET "sseg_sign[2]" IOSTANDARD = LVCMOS33;
NET "sseg_sign[1]" IOSTANDARD = LVCMOS33;
NET "sseg_sign[0]" IOSTANDARD = LVCMOS33;

# PlanAhead Generated physical constraints

NET "sseg_sign[6]" LOC = L18;
NET "sseg_sign[5]" LOC = T11;
NET "sseg_sign[4]" LOC = P15;
NET "sseg_sign[3]" LOC = K13;
NET "sseg_sign[2]" LOC = K16;
NET "sseg_sign[1]" LOC = R10;
NET "sseg_sign[0]" LOC = T10;

# PlanAhead Generated IO constraints

NET "clock" IOSTANDARD = LVCMOS33;
NET "kc" IOSTANDARD = LVCMOS33;
NET "kd" IOSTANDARD = LVCMOS33;
NET "reset" IOSTANDARD = LVCMOS33;

# PlanAhead Generated physical constraints

NET "clock" LOC = E3;
NET "kc" LOC = F4;
NET "kd" LOC = B2;
NET "reset" LOC = P18;
